//Ricky Gutierrez
//CSC137, Section 3
//Assignment #1
//mux4x1.v

module MuxMod(s0, s1, d0, d1, d2, d3, o);
	input s0, s1, d0, d1, d2, d3;
	output o;

	wire and0, and1, and2, and3;

	and(and0, ((~s0) & (~s1)), d0);
	and(and1, (s0 & (~s1)), d1);
	and(and2, ((~s0) & s1), d2);
	and(and3, (s0 & s1), d3);
	or(o, (and0 | and1), (and2 | and3));
endmodule

module TestMod;
	reg s0, s1, d0, d1, d2, d3;
	wire o;
	MuxMod my_mux(s0, s1, d0, d1, d2, d3, o);

	initial begin
		$display("Time\ts1\ts0\td0\td1\td2\td3\to");
		$display("---------------------------------------------------------");
		$monitor("%0d\t%b\t%b\t%b\t%b\t%b\t%b\t%b", $time, s1, s0, d0, d1, d2, d3, o);
	end

	initial begin
	//#1
		s0 = 0; s1 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 0; #1;
		s0 = 0; s1 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 1; #1;
		s0 = 0; s1 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 1; #1;
                s0 = 0; s1 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 0; #1;
                s0 = 0; s1 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 1; #1;
                s0 = 0; s1 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 1; #1;
	//#2
                s0 = 0; s1 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 1; #1;
                s0 = 0; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 1; #1;
                s0 = 0; s1 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 0; #1;
                s0 = 0; s1 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 1; #1;
                s0 = 0; s1 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 1; #1;
	//#3
		s0 = 1; s1 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 0; #1;
                s0 = 1; s1 = 0; d0 = 0; d1 = 0; d2 = 0; d3 = 1; #1;
                s0 = 1; s1 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 1; s1 = 0; d0 = 0; d1 = 0; d2 = 1; d3 = 1; #1;
                s0 = 1; s1 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 0; #1;
                s0 = 1; s1 = 0; d0 = 0; d1 = 1; d2 = 0; d3 = 1; #1;
                s0 = 1; s1 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 0; #1;
                s0 = 1; s1 = 0; d0 = 0; d1 = 1; d2 = 1; d3 = 1; #1;
	//#4
                s0 = 1; s1 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 0; #1;
                s0 = 1; s1 = 0; d0 = 1; d1 = 0; d2 = 0; d3 = 1; #1;
                s0 = 1; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 1; s1 = 0; d0 = 1; d1 = 0; d2 = 1; d3 = 1; #1;
                s0 = 1; s1 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 0; #1;
                s0 = 1; s1 = 0; d0 = 1; d1 = 1; d2 = 0; d3 = 1; #1;
                s0 = 1; s1 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 0; #1;
                s0 = 1; s1 = 0; d0 = 1; d1 = 1; d2 = 1; d3 = 1; #1;
	//#5
                s0 = 0; s1 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 0; #1;
                s0 = 0; s1 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 1; #1;
                s0 = 0; s1 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 1; #1;
                s0 = 0; s1 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 0; #1;
                s0 = 0; s1 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 1; #1;
                s0 = 0; s1 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 1; #1;
	//#6
		s0 = 0; s1 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 0; #1;
                s0 = 0; s1 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 1; #1;
                s0 = 0; s1 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 1; #1;
                s0 = 0; s1 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 0; #1;
                s0 = 0; s1 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 1; #1;
                s0 = 0; s1 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 0; #1;
                s0 = 0; s1 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 1; #1;
	//#7
                s0 = 1; s1 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 0; #1;
                s0 = 1; s1 = 1; d0 = 0; d1 = 0; d2 = 0; d3 = 1; #1;
                s0 = 1; s1 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 1; s1 = 1; d0 = 0; d1 = 0; d2 = 1; d3 = 1; #1;
                s0 = 1; s1 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 0; #1;
                s0 = 1; s1 = 1; d0 = 0; d1 = 1; d2 = 0; d3 = 1; #1;
                s0 = 1; s1 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 0; #1;
                s0 = 1; s1 = 1; d0 = 0; d1 = 1; d2 = 1; d3 = 1; #1;
	//#8
                s0 = 1; s1 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 0; #1;
                s0 = 1; s1 = 1; d0 = 1; d1 = 0; d2 = 0; d3 = 1; #1;
                s0 = 1; s1 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 0; #1;
                s0 = 1; s1 = 1; d0 = 1; d1 = 0; d2 = 1; d3 = 1; #1;
                s0 = 1; s1 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 0; #1;
                s0 = 1; s1 = 1; d0 = 1; d1 = 1; d2 = 0; d3 = 1; #1;
                s0 = 1; s1 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 0; #1;
                s0 = 1; s1 = 1; d0 = 1; d1 = 1; d2 = 1; d3 = 1; #1;
	end
endmodule
